-- COMPSYS 305 Miniproject
-- 2020 FPGPals
-- Modified by Cecil Symes, csym531

-- Displays text according to the current gamestate