library verilog;
use verilog.vl_types.all;
entity TextDisplay_vlg_vec_tst is
end TextDisplay_vlg_vec_tst;
