library verilog;
use verilog.vl_types.all;
entity TextDisplay_vlg_check_tst is
    port(
        pixel_on        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end TextDisplay_vlg_check_tst;
